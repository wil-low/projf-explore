`define CmdBranchTest          2  // BranchingTest
`define CmdFPGA         19  // FPGA routine
`define lblT7eq1         36  // Kill the Bit game: T7 == 1
`define CmdKillbits         51  // Kill the Bit game
`define CmdMaxSize        116  // Max file size
