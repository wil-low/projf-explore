// Infrared NEC protocol command codes
// full message: header, address, ~address, command, ~command

`define KEY_UP 8'h18
`define KEY_DOWN 8'h4A
`define KEY_LEFT 8'h10
`define KEY_RIGHT 8'h5A
`define KEY_OK 8'h38
`define KEY_1 8'hA2
`define KEY_2 8'h62
`define KEY_3 8'hE2
`define KEY_4 8'h22
`define KEY_5 8'h02
`define KEY_6 8'hC2
`define KEY_7 8'hE0
`define KEY_8 8'hA8
`define KEY_9 8'h90
`define KEY_0 8'h98
`define KEY_NUMERIC_STAR 8'h68
`define KEY_NUMERIC_POUND 8'hB0
