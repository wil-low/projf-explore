`define I_NOP0	4'b0000
`define I_LD	4'b0001
`define I_LDC	4'b0010
`define I_AND	4'b0011
`define I_ANDC	4'b0100
`define I_OR	4'b0101
`define I_ORC	4'b0110
`define I_XNOR	4'b0111
`define I_STO	4'b1000
`define I_STOC	4'b1001
`define I_IEN	4'b1010
`define I_OEN	4'b1011
`define I_JMP	4'b1100
`define I_RTN	4'b1101
`define I_SKZ	4'b1110
`define I_NOPF	4'b1111
