// Special circuit for LED drive control TM1638

`define TM1638_Display_Off 8'h80

`define TM1638_Display_1 8'h88
`define TM1638_Display_2 8'h89
`define TM1638_Display_3 8'h8a
`define TM1638_Display_4 8'h8b
`define TM1638_Display_5 8'h8c
`define TM1638_Display_6 8'h8d
`define TM1638_Display_7 8'h8e
`define TM1638_Display_8 8'h8f

`define TM1638_AutoIncrementMode 8'h40

`define TM1638_SetAddress 8'hc0
