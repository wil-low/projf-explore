`define CCHAR0 8'h80
`define CCHAR1 8'h81
`define CCHAR2 8'h82
`define CCHAR3 8'h83
`define CCHAR4 8'h84
`define CCHAR5 8'h85
`define CCHAR6 8'h86
`define CCHAR7 8'h87
